// This file (bs_smoke_test.sv) will be included within bs_test_pkg.sv.
// It assumes barrel_shifter_base_test, bs_env, and bs_random_stimulus_sequence types
// are available via prior includes in the package.

class bs_smoke_test extends barrel_shifter_base_test;
  `uvm_component_utils(bs_smoke_test)

  // Environment handle.
  // The parameters used for declaration (32, 1) must match the parameters
  // used during actual instantiation, which are derived from cfg_dut_data_width
  // and cfg_effective_latency after super.build_phase().
  // This test ensures they match by setting them via uvm_config_db before super.build_phase().
  bs_env #(32, 1) env_h; // DATA_WIDTH=32, Effective Latency=1 (derived from NUM_STAGES=1)

  function new(string name = "bs_smoke_test", uvm_component parent = null);
    super.new(name, parent);
  endfunction

  virtual function void build_phase(uvm_phase phase);
    `uvm_info(get_type_name(), "Build phase of smoke test", UVM_MEDIUM)
    // Set the desired configuration for this specific test.
    // These values will be read by barrel_shifter_base_test's build_phase.
    // This ensures this test runs with DATA_WIDTH=32 and NUM_STAGES=1 (effective latency 1).
    uvm_config_db#(int)::set(this, "", "dut_data_width", 32);
    uvm_config_db#(int)::set(this, "", "dut_num_stages", 1); // This results in cfg_effective_latency = 1

    // Call base class's build_phase to read these configurations (and others)
    // and calculate cfg_dut_data_width and cfg_effective_latency.
    super.build_phase(phase); 
    // Now, cfg_dut_data_width in the base class is 32.
    // And cfg_effective_latency in the base class is 1 (since cfg_dut_num_stages was set to 1).

    // Create the environment, parameterized with the values determined by the base class build.
    // The type of env_h (bs_env#(32,1)) must be compatible with these parameters.
    // Since cfg_dut_data_width is 32 and cfg_effective_latency is 1, this is consistent.
    env_h = bs_env#(cfg_dut_data_width, cfg_effective_latency)::type_id::create("env", this);
    if (env_h == null) begin
      `uvm_fatal(get_type_name(), "Environment creation failed in smoke test.")
    end
    // Optional: if base class had a generic handle like `super.env_inst` for uvm_env
    // super.env_inst = env_h; 
  endfunction

  virtual task run_phase(uvm_phase phase);
    // Sequence handle, parameterized by the DATA_WIDTH of the environment instance.
    bs_random_stimulus_sequence#(env_h.DATA_WIDTH) seq; 
    
    phase.raise_objection(this, "Smoke test starting");
    `uvm_info(get_type_name(), "Smoke test run_phase starting", UVM_MEDIUM)

    // Create the sequence instance
    seq = bs_random_stimulus_sequence#(env_h.DATA_WIDTH)::type_id::create("seq");
    if (seq == null) begin
       `uvm_fatal(get_type_name(), "Sequence creation failed")
    end

    seq.num_transactions = 5; // Smoke test runs a few transactions
    
    // Start the sequence on the agent's sequencer via the env handle
    if (env_h == null || env_h.agent == null || env_h.agent.sequencer == null) begin
      `uvm_fatal(get_type_name(), "Environment, agent, or sequencer handle is null. Cannot start sequence.")
    end
    seq.start(env_h.agent.sequencer);
    
    // A small delay to allow sequence to complete and items to drain through scoreboard.
    // UVM objections raised by the sequence (via start_item/finish_item) and driver
    // should ideally manage the simulation end time correctly.
    // This extra delay is a safety net, can be very small or removed if objections are robust.
    #200ns; 
    
    `uvm_info(get_type_name(), "Smoke test run_phase finishing", UVM_MEDIUM)
    phase.drop_objection(this, "Smoke test finished");
  endtask

endclass
