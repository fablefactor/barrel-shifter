// This file (bs_full_rotate_sequence.sv) will be included within bs_test_pkg.sv.

class bs_full_rotate_sequence #(
  parameter DATA_WIDTH = 32
) extends uvm_sequence #(bs_transaction#(DATA_WIDTH));

  `uvm_object_param_utils(bs_full_rotate_sequence#(DATA_WIDTH))

  int num_transactions = 10; 

  function new(string name = "bs_full_rotate_sequence");
    super.new(name);
  endfunction

  virtual task body();
    bs_transaction#(DATA_WIDTH) m_req;
    
    if (num_transactions <= 0) begin
      `uvm_warning(get_type_name(), $sformatf("num_transactions is %0d, sequence will not send any items.", num_transactions))
      return;
    end

    `uvm_info(get_type_name(), $sformatf("Starting full_rotate_sequence: generating %0d transactions (shift_amount=0).", num_transactions), UVM_MEDIUM)

    for (int i = 0; i < num_transactions; i++) begin
      `uvm_create(m_req)
      start_item(m_req);
      // A "full rotate" where data returns to original position means shift_amount is 0 
      // or a multiple of DATA_WIDTH. Given shift_amount width is $clog2(DATA_WIDTH) (or 1 if DATA_WIDTH=1),
      // and the transaction constraint `shift_amount < DATA_WIDTH`,
      // only 0 is consistently representable and valid for this behavior across all DATA_WIDTH.
      if (!m_req.randomize() with { shift_amount == '0; }) begin 
        `uvm_error(get_type_name(), "Failed to randomize transaction with shift_amount == 0 for full_rotate_sequence")
      end else begin
        `uvm_info(get_type_name(), $sformatf("Sent full_rotate transaction %0d/%0d: %s", i+1, num_transactions, m_req.convert2string()), UVM_HIGH)
      end
      finish_item(m_req);
    end
    `uvm_info(get_type_name(), $sformatf("Finished full_rotate_sequence after %0d transactions.", num_transactions), UVM_MEDIUM)
  endtask

endclass
