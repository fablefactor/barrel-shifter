// This file (base_test.sv) will be included within bs_test_pkg.sv,
// so uvm_pkg import and uvm_macros.svh include are via the package.
// It assumes bs_env type is available via prior include in the package.

class barrel_shifter_base_test extends uvm_test;
  `uvm_component_utils(barrel_shifter_base_test)

  // Configuration values read from uvm_config_db, with defaults
  protected int cfg_dut_data_width = 32;
  protected int cfg_dut_num_stages = 1;   // This is the NUM_STAGES parameter of the DUT itself
  protected int cfg_effective_latency = 1; // Monitor latency: max(1, cfg_dut_num_stages)

  function new(string name = "barrel_shifter_base_test", uvm_component parent = null);
    super.new(name, parent);
  endfunction

  virtual function void build_phase(uvm_phase phase);
    string current_test_name = get_full_name(); // For more specific logging messages
    super.build_phase(phase);

    // Get DATA_WIDTH for the DUT
    if (!uvm_config_db#(int)::get(this, "", "dut_data_width", cfg_dut_data_width)) begin
      `uvm_info(get_type_name(), $sformatf("[%s] 'dut_data_width' not set via uvm_config_db. Using default: %0d.", current_test_name, cfg_dut_data_width), UVM_MEDIUM)
    end

    // Get NUM_STAGES for the DUT (the Verilog module parameter)
    if (!uvm_config_db#(int)::get(this, "", "dut_num_stages", cfg_dut_num_stages)) begin
      `uvm_info(get_type_name(), $sformatf("[%s] 'dut_num_stages' not set via uvm_config_db. Using default: %0d.", current_test_name, cfg_dut_num_stages), UVM_MEDIUM)
    end

    // Validate dut_data_width
    if (cfg_dut_data_width <= 0) begin
      `uvm_fatal(get_type_name(), $sformatf("[%s] Configured 'dut_data_width' (%0d) must be greater than 0.", current_test_name, cfg_dut_data_width))
    end
    
    // dut_num_stages from DUT Verilog can be 0 (treated as 1 stage/cycle latency by DUT).
    // Calculate effective latency for the monitor based on DUT's NUM_STAGES parameter.
    // If DUT NUM_STAGES is 0, effective latency is 1. Otherwise, it's NUM_STAGES.
    // This interpretation should match how barrel_shifter.v handles NUM_STAGES = 0.
    cfg_effective_latency = (cfg_dut_num_stages == 0) ? 1 : cfg_dut_num_stages;
    // An alternative, if cfg_dut_num_stages could be negative or uninitialized from Verilog side:
    // cfg_effective_latency = (cfg_dut_num_stages <= 0) ? 1 : cfg_dut_num_stages;
    // Given Verilog parameter constraints, NUM_STAGES>=0 is expected.

    `uvm_info(get_type_name(), 
              $sformatf("[%s] Test Configuration: DUT_DATA_WIDTH=%0d, DUT_NUM_STAGES_PARAM=%0d, Effective Monitor Latency=%0d.",
                        current_test_name, cfg_dut_data_width, cfg_dut_num_stages, cfg_effective_latency), UVM_LOW);
    
    // Derived tests will use cfg_dut_data_width and cfg_effective_latency 
    // to instantiate a bs_env#(cfg_dut_data_width, cfg_effective_latency).
    // They will also set these parameters into the uvm_config_db for the env to pick up
    // if the env itself needs them for some reason (though bs_env uses its own parameters).
  endfunction

  // Default run_phase. Derived tests will typically start sequences here.
  virtual task run_phase(uvm_phase phase);
    phase.raise_objection(this, {get_full_name(), " base test starting now"});
    // A minimal delay to keep simulation alive if no sequences are run by derived tests
    // or if derived test forgets to call super.run_phase() but doesn't implement its own objection.
    #100ns; 
    phase.drop_objection(this, {get_full_name(), " base test finishing now"});
  endtask

  virtual function void end_of_elaboration_phase(uvm_phase phase);
    super.end_of_elaboration_phase(phase);
    `uvm_info(get_type_name(), $sformatf("[%s] Printing UVM topology...", get_full_name()), UVM_LOW);
    uvm_top.print_topology();
  endfunction

endclass
